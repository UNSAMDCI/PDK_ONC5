* HSPICE netlist generated with ICnet by 'unsam' on Mon Oct 24 2016 at 10:32:55

*
* MAIN CELL: Component pathname : $BASIC_CELLS_ONC5/D_CELLS/AND3X1
*
.subckt AND3X1  D_GND D_VDD OUT A B C

        M_ENM2 N_17_ESC1 B N_19_ESC2 D_GND enm w=2.4u l=0.6u m=1 mult=1 region=1
        M_ENM1 N_24_ESC3 A N_17_ESC1 D_GND enm w=2.4u l=0.6u m=1 mult=1 region=1
        M_EPM2 N_24_ESC3 A D_VDD D_VDD epm w=2.4u l=0.6u m=1 mult=1 region=1
        M_EPM1 N_24_ESC3 B D_VDD D_VDD epm w=2.4u l=0.6u m=1 mult=1 region=1
        M_ENM4 OUT N_24_ESC3 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 region=1
        M_EPM4 OUT N_24_ESC3 D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 region=1
        M_ENM3 N_19_ESC2 C D_GND D_GND enm w=2.4u l=0.6u m=1 mult=1 region=1
        M_EPM3 N_24_ESC3 C D_VDD D_VDD epm w=2.4u l=0.6u m=1 mult=1 region=1
.ends AND3X1

