* HSPICE netlist generated with ICnet by 'unsam' on Wed Feb  1 2017 at 09:14:41

*
* MAIN CELL: Component pathname : $BASIC_CELLS_ONC5/D_CELLS/BUX4
*
.subckt BUX4  D_GND D_VDD OUT IN

        M_EPM2 OUT N_2_ESC1 D_VDD D_VDD epm w=2.75u l=0.6u m=7 mult=7 
        M_ENM2 OUT N_2_ESC1 D_GND D_GND enm w=1.6u l=0.6u m=6 mult=6 
        M_EPM1 N_2_ESC1 IN D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1
        M_ENM1 N_2_ESC1 IN D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
.ends BUX4

