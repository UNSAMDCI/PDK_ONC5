* HSPICE netlist generated with ICnet by 'unsam' on Fri Mar 31 2017 at 08:51:37

*
* MAIN CELL: Component pathname : $BASIC_CELLS_ONC5/D_CELLS/NO4X1
*
.subckt NO4X1  OUT A B C D D_GND D_VDD

        M_EPM7 OUT OR D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_ENM7 OUT OR D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM6 N_74_ESC1 OUT2 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM5 OR OUT1 N_74_ESC1 D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM6 OR OUT2 D_VDD D_VDD epm w=0.8u l=0.6u m=1 mult=1 
        M_EPM5 OR OUT1 D_VDD D_VDD epm w=0.8u l=0.6u m=1 mult=1 
        M_ENM4 OUT2 D D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM3 OUT2 C D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM4 N_25_ESC2 C D_VDD D_VDD epm w=3.2u l=0.6u m=1 mult=1 
        M_EPM3 OUT2 D N_25_ESC2 D_VDD epm w=3.2u l=0.6u m=1 mult=1 
        M_ENM2 OUT1 B D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM1 OUT1 A D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM2 N_14_ESC3 A D_VDD D_VDD epm w=3.2u l=0.6u m=1 mult=1 
        M_EPM1 OUT1 B N_14_ESC3 D_VDD epm w=3.2u l=0.6u m=1 mult=1 
.ends NO4X1

