* LVS netlist generated with ICnet by 'unsam' on Wed Jan 25 2017 at 12:35:40

*
* Component pathname : $BASIC_CELLS_ONC5/D_CELLS/GATES/inv
*
.subckt inv  OUT D_GND D_VDD IN

        M_ENM1 OUT IN D_GND D_GND enm m=1 W=0.8u L=0.6u
        M_EPM1 OUT IN D_VDD D_VDD epm m=1 W=1.6u L=0.6u
.ends inv

*
* Component pathname : $BASIC_CELLS_ONC5/D_CELLS/FAX1
*
.subckt FAX1  CO S D_GND D_VDD A B CI

        M_I$25 N$89 B D_GND D_GND enm m=1 W=0.8u L=0.6u
        M_I$24 N$102 N$16 N$89 D_GND enm m=1 W=0.8u L=0.6u
        M_I$23 N$89 CI D_GND D_GND enm m=1 W=0.8u L=0.6u
        X_INV2 CO D_GND D_VDD N$16 inv
        X_INV1 S D_GND D_VDD N$102 inv
        M_I$29 N$102 CI N$84 D_GND enm m=1 W=0.8u L=0.6u
        M_I$19 N$80 B N$76 D_VDD epm m=1 W=1.6u L=0.6u
        M_I$18 N$76 A D_VDD D_VDD epm m=1 W=1.6u L=0.6u
        M_I$17 N$65 A D_VDD D_VDD epm m=1 W=1.6u L=0.6u
        M_I$16 N$102 N$16 N$65 D_VDD epm m=1 W=1.6u L=0.6u
        M_I$15 N$65 B D_VDD D_VDD epm m=1 W=1.6u L=0.6u
        M_I$14 N$65 CI D_VDD D_VDD epm m=1 W=1.6u L=0.6u
        M_I$10 N$3 A D_GND D_GND enm m=1 W=0.8u L=0.6u
        M_I$9 N$3 B D_GND D_GND enm m=1 W=0.8u L=0.6u
        M_I$8 N$16 CI N$3 D_GND enm m=1 W=0.8u L=0.6u
        M_I$7 N$14 A D_GND D_GND enm m=1 W=0.8u L=0.6u
        M_I$6 N$16 B N$14 D_GND enm m=1 W=0.8u L=0.6u
        M_I$5 N$20 A D_VDD D_VDD epm m=1 W=1.6u L=0.6u
        M_I$4 N$20 B D_VDD D_VDD epm m=1 W=1.6u L=0.6u
        M_I$3 N$16 CI N$20 D_VDD epm m=1 W=1.6u L=0.6u
        M_I$2 N$16 B N$32 D_VDD epm m=1 W=1.6u L=0.6u
        M_I$1 N$32 A D_VDD D_VDD epm m=1 W=1.6u L=0.6u
        M_I$20 N$102 CI N$80 D_VDD epm m=1 W=1.6u L=0.6u
        M_I$28 N$84 B N$57 D_GND enm m=1 W=0.8u L=0.6u
        M_I$27 N$57 A D_GND D_GND enm m=1 W=0.8u L=0.6u
        M_I$26 N$89 A D_GND D_GND enm m=1 W=0.8u L=0.6u
.ends FAX1

