* HSPICE netlist generated with ICnet by 'unsam' on Fri Mar 31 2017 at 08:56:28

*
* MAIN CELL: Component pathname : $BASIC_CELLS_ONC5/D_CELLS/NO6X1
*
.subckt NO6X1  OUT A B C D D_GND D_VDD E F

        M_ENM9 OUT2 F D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM9 OUT2 F N_90_ESC1 D_VDD epm w=4.5u l=0.6u m=1 mult=1 
        M_ENM8 OUT1 E D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM8 OUT1 E N_77_ESC2 D_VDD epm w=4.5u l=0.6u m=1 mult=1 
        M_EPM7 OUT OR D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_ENM7 OUT OR D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM6 N_74_ESC3 OUT2 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM5 OR OUT1 N_74_ESC3 D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM6 OR OUT2 D_VDD D_VDD epm w=0.8u l=0.6u m=1 mult=1 
        M_EPM5 OR OUT1 D_VDD D_VDD epm w=0.8u l=0.6u m=1 mult=1 
        M_ENM4 OUT2 D D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM3 OUT2 C D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM4 N_25_ESC4 C D_VDD D_VDD epm w=4.5u l=0.6u m=1 mult=1 
        M_EPM3 N_90_ESC1 D N_25_ESC4 D_VDD epm w=4.5u l=0.6u m=1 mult=1 
        M_ENM2 OUT1 B D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM1 OUT1 A D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM2 N_14_ESC5 A D_VDD D_VDD epm w=4.5u l=0.6u m=1 mult=1 
        M_EPM1 N_77_ESC2 B N_14_ESC5 D_VDD epm w=4.5u l=0.6u m=1 mult=1 
.ends NO6X1

