* HSPICE netlist generated with ICnet by 'unsam' on Mon Oct 24 2016 at 10:39:20

*
* MAIN CELL: Component pathname : $BASIC_CELLS_ONC5/D_CELLS/AO222X1
*
.subckt AO222X1  D_GND D_VDD OUT A B C D E F

        M_ENM12 N_61_ESC1 OR3 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM11 N_61_ESC1 OR2 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM10 N_61_ESC1 OR1 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM12 N_61_ESC1 OR3 N_29_ESC2 D_VDD epm w=4.8u l=0.6u m=1 mult=1
        M_EPM11 N_29_ESC2 OR2 N_31_ESC3 D_VDD epm w=4.8u l=0.6u m=1 mult=1
        M_EPM10 N_31_ESC3 OR1 D_VDD D_VDD epm w=4.8u l=0.6u m=1 mult=1 
        M_EPM9 OR3 N_20_ESC4 D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_ENM9 OR3 N_20_ESC4 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM8 N_25_ESC5 F D_GND D_GND enm w=1.6u l=0.6u m=1 mult=1
        M_ENM7 N_20_ESC4 E N_25_ESC5 D_GND enm w=1.6u l=0.6u m=1 mult=1 
        M_EPM8 N_20_ESC4 E D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_EPM7 N_20_ESC4 F D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_ENM6 OR2 N_11_ESC6 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM5 N_16_ESC7 D D_GND D_GND enm w=1.6u l=0.6u m=1 mult=1 
        M_ENM4 N_11_ESC6 C N_16_ESC7 D_GND enm w=1.6u l=0.6u m=1 mult=1 
        M_EPM5 N_11_ESC6 C D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_EPM4 N_11_ESC6 D D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_EPM3 OR1 N_2_ESC8 D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_ENM3 OR1 N_2_ESC8 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM6 OR2 N_11_ESC6 D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_ENM2 N_7_ESC9 B D_GND D_GND enm w=1.6u l=0.6u m=1 mult=1 
        M_ENM1 N_2_ESC8 A N_7_ESC9 D_GND enm w=1.6u l=0.6u m=1 mult=1
        M_EPM2 N_2_ESC8 A D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_EPM1 N_2_ESC8 B D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_EPM13 OUT N_61_ESC1 D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_ENM13 OUT N_61_ESC1 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
.ends AO222X1

