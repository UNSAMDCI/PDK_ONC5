* HSPICE netlist generated with ICnet by 'unsam' on Mon Oct 24 2016 at 10:49:26

*
* MAIN CELL: Component pathname : $BASIC_CELLS_ONC5/D_CELLS/OA211X1
*
.subckt OA211X1  D_GND D_VDD OUT A B C D

        M_EPM7 OR_O N_27_ESC1 D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 region=1
        M_ENM7 OR_O N_27_ESC1 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 region=1
        M_ENM6 N_27_ESC1 B D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 region=1
        M_ENM5 N_27_ESC1 A D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 region=1
        M_EPM6 N_29_ESC2 A D_VDD D_VDD epm w=3.2u l=0.6u m=1 mult=1 region=1
        M_EPM5 N_27_ESC1 B N_29_ESC2 D_VDD epm w=3.2u l=0.6u m=1 mult=1 region=1
        M_ENM1 N_2_ESC3 OR_O N_7_ESC4 D_GND enm w=2.4u l=0.6u m=1 mult=1 region=1
        M_ENM4 OUT N_2_ESC3 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 region=1
        M_EPM3 N_2_ESC3 C D_VDD D_VDD epm w=2.4u l=0.6u m=1 mult=1 region=1
        M_ENM3 N_9_ESC5 C D_GND D_GND enm w=2.4u l=0.6u m=1 mult=1 region=1
        M_ENM2 N_7_ESC4 D N_9_ESC5 D_GND enm w=2.4u l=0.6u m=1 mult=1 region=1
        M_EPM4 OUT N_2_ESC3 D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 region=1
        M_EPM2 N_2_ESC3 OR_O D_VDD D_VDD epm w=2.4u l=0.6u m=1 mult=1 region=1
        M_EPM1 N_2_ESC3 D D_VDD D_VDD epm w=2.4u l=0.6u m=1 mult=1 region=1
.ends OA211X1

