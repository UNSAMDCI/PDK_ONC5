* HSPICE netlist generated with ICnet by 'unsam' on Mon Oct 24 2016 at 10:47:01

*
* MAIN CELL: Component pathname : $BASIC_CELLS_ONC5/D_CELLS/NA3I1X1

.subckt NA3I1X1  D_GND D_VDD OUT B C NA

        M_EPM4 A NA D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 region=1
        M_EPM3 OUT C D_VDD D_VDD epm w=2.4u l=0.6u m=1 mult=1 region=1
        M_ENM3 N_9_ESC1 C D_GND D_GND enm w=2.4u l=0.6u m=1 mult=1 region=1
        M_ENM4 A NA D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 region=1 
        M_ENM2 N_7_ESC2 B N_9_ESC1 D_GND enm w=2.4u l=0.6u m=1 mult=1 region=1
        M_ENM1 OUT A N_7_ESC2 D_GND enm w=2.4u l=0.6u m=1 mult=1 region=1
        M_EPM2 OUT A D_VDD D_VDD epm w=2.4u l=0.6u m=1 mult=1 region=1
        M_EPM1 OUT B D_VDD D_VDD epm w=2.4u l=0.6u m=1 mult=1 region=1 
.ends NA3I1X1

