* HSPICE netlist generated with ICnet by 'unsam' on Fri Mar 31 2017 at 08:58:19

*
* MAIN CELL: Component pathname : $BASIC_CELLS_ONC5/D_CELLS/OR2x1
*
.subckt OR2X1  D_GND D_VDD OUT A B

        M_ENM3 OUT NOOUT D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM3 OUT NOOUT D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_ENM2 NOOUT B D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM1 NOOUT A D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM2 N_14_ESC1 A D_VDD D_VDD epm w=3.2u l=0.6u m=1 mult=1 
        M_EPM1 NOOUT B N_14_ESC1 D_VDD epm w=3.2u l=0.6u m=1 mult=1 
.ends OR2X1

