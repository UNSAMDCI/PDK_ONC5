* HSPICE netlist generated with ICnet by 'unsam' on Wed Feb  1 2017 at 12:10:37

*
* MAIN CELL: Component pathname : $BASIC_CELLS_ONC5/D_CELLS/BUX8
*
.subckt BUX8  D_GND D_VDD Z IN

        M_EPM2 Z N_2_ESC1 D_VDD D_VDD epm w=38.4u l=0.6u m=1 mult=1 
        M_ENM2 Z N_2_ESC1 D_GND D_GND enm w=19.2u l=0.6u m=1 mult=1 
        M_EPM1 N_2_ESC1 IN D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_ENM1 N_2_ESC1 IN D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
.ends BUX8

