* HSPICE netlist generated with ICnet by 'unsam' on Mon Oct 24 2016 at 10:44:53

*
* MAIN CELL: Component pathname : $BASIC_CELLS_ONC5/D_CELLS/AO32X1
*
.subckt AO32X1  D_GND D_VDD OUT A B C D E

        M_EPM10 OUT N_27_ESC1 D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 region=1
        M_ENM10 OUT N_27_ESC1 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 region=1
        M_ENM9 N_27_ESC1 AND_O2 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 region=1
        M_ENM8 N_27_ESC1 AND_O1 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 region=1
        M_EPM9 N_29_ESC2 AND_O1 D_VDD D_VDD epm w=3.2u l=0.6u m=1 mult=1 region=1
        M_EPM8 N_27_ESC1 AND_O2 N_29_ESC2 D_VDD epm w=3.2u l=0.6u m=1 mult=1
        M_ENM7 AND_O2 N_17_ESC3 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 region=1
        M_ENM6 N_22_ESC4 E D_GND D_GND enm w=1.6u l=0.6u m=1 mult=1 region=1
        M_ENM5 N_17_ESC3 D N_22_ESC4 D_GND enm w=1.6u l=0.6u m=1 mult=1 region=1
        M_EPM6 N_17_ESC3 D D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 region=1
        M_EPM5 N_17_ESC3 E D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 region=1
        M_EPM7 AND_O2 N_17_ESC3 D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 region=1
        M_EPM4 AND_O1 N_2_ESC5 D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 region=1
        M_ENM4 AND_O1 N_2_ESC5 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 region=1
        M_EPM3 N_2_ESC5 C D_VDD D_VDD epm w=2.4u l=0.6u m=1 mult=1 region=1
        M_ENM3 N_9_ESC6 C D_GND D_GND enm w=2.4u l=0.6u m=1 mult=1 region=1
        M_ENM2 N_7_ESC7 B N_9_ESC6 D_GND enm w=2.4u l=0.6u m=1 mult=1 region=1
        M_ENM1 N_2_ESC5 A N_7_ESC7 D_GND enm w=2.4u l=0.6u m=1 mult=1 region=1
        M_EPM2 N_2_ESC5 A D_VDD D_VDD epm w=2.4u l=0.6u m=1 mult=1 region=1
        M_EPM1 N_2_ESC5 B D_VDD D_VDD epm w=2.4u l=0.6u m=1 mult=1 region=1
.ends AO32X1

