* HSPICE netlist generated with ICnet by 'unsam' on Fri Mar 31 2017 at 08:44:04

*
* MAIN CELL: Component pathname : $BASIC_CELLS_ONC5/D_CELLS/NA4X1
*
.subckt NA4X1  OUT A B C D D_GND D_VDD

        M_ENM7 OUT N_108_ESC1 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM4 OUT2 C D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_EPM3 OUT2 D D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_ENM3 N_106_ESC2 B D_GND D_GND enm w=1.6u l=0.6u m=1 mult=1 
        M_ENM1 OUT1 A N_106_ESC2 D_GND enm w=1.6u l=0.6u m=1 mult=1 
        M_EPM2 OUT1 A D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_EPM1 OUT1 B D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_EPM7 OUT N_108_ESC1 D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_EPM5 N_108_ESC1 OUT2 N_122_ESC3 D_VDD epm w=6.4u l=0.6u m=1 mult=1
        M_ENM6 N_108_ESC1 OUT2 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM4 N_115_ESC4 D D_GND D_GND enm w=1.6u l=0.6u m=1 mult=1 
        M_ENM2 OUT2 C N_115_ESC4 D_GND enm w=1.6u l=0.6u m=1 mult=1 
        M_ENM5 N_108_ESC1 OUT1 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM6 N_122_ESC3 OUT1 D_VDD D_VDD epm w=6.4u l=0.6u m=1 mult=1 
.ends NA4X1

