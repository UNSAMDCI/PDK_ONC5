* HSPICE netlist generated with ICnet by 'unsam' on Wed Nov 16 2016 at 08:49:18

*
* Component pathname : $BASIC_CELLS_ONC5/D_CELLS/MU2IX1
*
.subckt MU2IX1  QN D_GND D_VDD IN0 IN1 S

        M_EPM5 CLK1 S D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_ENM5 CLK1 S D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1  
        M_EPM4 N_25_ESC1 IN1 D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_EPM3 QN CLK1 N_25_ESC1 D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_ENM4 N_21_ESC2 IN1 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM3 QN S N_21_ESC2 D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM2 N_2_ESC3 IN0 D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_EPM1 QN S N_2_ESC3 D_VDD epm w=1.6u l=0.6u m=1 mult=1 
        M_ENM2 N_6_ESC4 IN0 D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_ENM1 QN CLK1 N_6_ESC4 D_GND enm w=0.8u l=0.6u m=1 mult=1 
.ends MU2IX1

