* HSPICE netlist generated with ICnet by 'unsam' on Wed Feb  1 2017 at 11:40:51

*
* MAIN CELL: Component pathname : $BASIC_CELLS_ONC5/D_CELLS/DLY1p6LX1
*
.subckt DLY1P6LX1  Q D_GND D_VDD D

        M_ENM3 Q N_146_ESC1 D_GND D_GND enm w=2.4u l=0.6u m=1 mult=1 
        M_EPM4 Q N_146_ESC1 D_VDD D_VDD epm w=4.8u l=0.6u m=1 mult=1 
        M_ENM2 N_146_ESC1 N_147_ESC2 D_GND D_GND enm w=1.4u l=1.55u m=1 mult=1
        M_EPM2 N_146_ESC1 N_147_ESC2 D_VDD D_VDD epm w=3.4u l=1.55u m=1 mult=1
        M_ENM1 N_147_ESC2 N_7_ESC3 D_GND D_GND enm w=1.4u l=1.55u m=1 mult=1
        M_EPM1 N_147_ESC2 N_7_ESC3 D_VDD D_VDD epm w=3.4u l=1.55u m=1 mult=1
        M_ENM7 N_7_ESC3 D D_GND D_GND enm w=0.8u l=0.6u m=1 mult=1 
        M_EPM3 N_7_ESC3 D D_VDD D_VDD epm w=1.6u l=0.6u m=1 mult=1 
.ends DLY1P6LX1

